// $Id: $
// File name:   sensor_s.sv
// Created:     1/21/2020
// Author:      Haoming Duan
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: This file is a structural coding of sensor error detector, which has two ports, input sensors[3:0] and output error
